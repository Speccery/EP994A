----------------------------------------------------------------------------------
-- Engineer:	Erik Piehl 
-- 
-- Create Date:    07:01:30 04/15/2017 
-- Design Name: 	 testrom.vhd
-- Module Name:    testrom - Behavioral 
-- Project Name: 	 TMS9900 Test ROM code
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity testrom is
    Port ( clk : in  STD_LOGIC;
           addr : in  STD_LOGIC_VECTOR (7 downto 0);
           data_out : out  STD_LOGIC_VECTOR (15 downto 0));
end testrom;

architecture Behavioral of testrom is
	constant romLast : integer := 4095;
	type pgmRomArray is array(0 to romLast) of STD_LOGIC_VECTOR (15 downto 0);
	constant pgmRom : pgmRomArray := (  
            x"8300"
           ,x"0046"
           ,x"a000"
           ,x"0020"
           ,x"a000"
           ,x"0020"
           ,x"8320"
           ,x"046a"
           ,x"8320"
           ,x"0458"
           ,x"8320"
           ,x"049c"
           ,x"8320"
           ,x"04ac"
           ,x"8340"
           ,x"04da"
           ,x"0300"
           ,x"0000"
           ,x"0580"
           ,x"04cc"
           ,x"3402"
           ,x"1f02"
           ,x"1603"
           ,x"0203"
           ,x"ffff"
           ,x"1002"
           ,x"0203"
           ,x"1234"
           ,x"d060"
           ,x"8802"
           ,x"0205"
           ,x"0100"
           ,x"b805"
           ,x"8379"
           ,x"0380"
           ,x"0300"
           ,x"0000"
           ,x"02e0"
           ,x"8300"
           ,x"04e0"
           ,x"a000"
           ,x"d803"
           ,x"8c00"
           ,x"0201"
           ,x"051c"
           ,x"0202"
           ,x"8000"
           ,x"d831"
           ,x"8c02"
           ,x"d802"
           ,x"8c02"
           ,x"0222"
           ,x"0100"
           ,x"0282"
           ,x"8800"
           ,x"16f7"
           ,x"04c0"
           ,x"0201"
           ,x"4000"
           ,x"06c1"
           ,x"d801"
           ,x"8c02"
           ,x"06c1"
           ,x"d801"
           ,x"8c02"
           ,x"d800"
           ,x"8c00"
           ,x"0601"
           ,x"16fc"
           ,x"06a0"
           ,x"03f2"
           ,x"0200"
           ,x"0380"
           ,x"06a0"
           ,x"038a"
           ,x"0201"
           ,x"0020"
           ,x"0202"
           ,x"1700"
           ,x"d802"
           ,x"8c00"
           ,x"0601"
           ,x"16fc"
           ,x"1028"
           ,x"04e0"
           ,x"8320"
           ,x"04c1"
           ,x"0202"
           ,x"1234"
           ,x"0203"
           ,x"ffff"
           ,x"0204"
           ,x"2000"
           ,x"0205"
           ,x"0014"
           ,x"0206"
           ,x"def0"
           ,x"0207"
           ,x"3300"
           ,x"c801"
           ,x"8322"
           ,x"0420"
           ,x"0010"
           ,x"d804"
           ,x"8322"
           ,x"0420"
           ,x"0014"
           ,x"c181"
           ,x"0586"
           ,x"d807"
           ,x"8322"
           ,x"0420"
           ,x"0014"
           ,x"0606"
           ,x"16fa"
           ,x"0420"
           ,x"000c"
           ,x"0524"
           ,x"0581"
           ,x"0241"
           ,x"001f"
           ,x"0281"
           ,x"0018"
           ,x"16e7"
           ,x"0200"
           ,x"0040"
           ,x"c800"
           ,x"8320"
           ,x"0200"
           ,x"1234"
           ,x"0209"
           ,x"0003"
           ,x"0420"
           ,x"000c"
           ,x"1912"
           ,x"d800"
           ,x"9c02"
           ,x"06c0"
           ,x"d800"
           ,x"9c02"
           ,x"06c0"
           ,x"04c1"
           ,x"d060"
           ,x"9800"
           ,x"d0a0"
           ,x"9800"
           ,x"0982"
           ,x"e042"
           ,x"c801"
           ,x"8322"
           ,x"0420"
           ,x"0010"
           ,x"04c1"
           ,x"d060"
           ,x"9800"
           ,x"d0a0"
           ,x"9800"
           ,x"0982"
           ,x"e042"
           ,x"c801"
           ,x"8322"
           ,x"0420"
           ,x"0010"
           ,x"04c1"
           ,x"d060"
           ,x"9802"
           ,x"d0a0"
           ,x"9802"
           ,x"0982"
           ,x"e042"
           ,x"c801"
           ,x"8322"
           ,x"0420"
           ,x"0010"
           ,x"0220"
           ,x"2000"
           ,x"0609"
           ,x"16d2"
           ,x"04cc"
           ,x"1e00"
           ,x"1d02"
           ,x"0300"
           ,x"0002"
           ,x"0203"
           ,x"03e8"
           ,x"04c0"
           ,x"c800"
           ,x"8320"
           ,x"020c"
           ,x"0024"
           ,x"30c0"
           ,x"020c"
           ,x"0006"
           ,x"3601"
           ,x"c801"
           ,x"8322"
           ,x"0420"
           ,x"0010"
           ,x"0420"
           ,x"000c"
           ,x"0524"
           ,x"0220"
           ,x"0100"
           ,x"0280"
           ,x"0600"
           ,x"16ee"
           ,x"c060"
           ,x"a000"
           ,x"c801"
           ,x"8322"
           ,x"0420"
           ,x"0010"
           ,x"0420"
           ,x"000c"
           ,x"0524"
           ,x"0420"
           ,x"000c"
           ,x"1905"
           ,x"c060"
           ,x"a004"
           ,x"c801"
           ,x"8322"
           ,x"0420"
           ,x"0010"
           ,x"0420"
           ,x"000c"
           ,x"0524"
           ,x"c060"
           ,x"a006"
           ,x"c801"
           ,x"8322"
           ,x"0420"
           ,x"0010"
           ,x"0420"
           ,x"000c"
           ,x"0524"
           ,x"04cc"
           ,x"3401"
           ,x"c801"
           ,x"8322"
           ,x"0420"
           ,x"0010"
           ,x"0420"
           ,x"000c"
           ,x"0524"
           ,x"0603"
           ,x"16c2"
           ,x"c060"
           ,x"6000"
           ,x"0281"
           ,x"aa01"
           ,x"1607"
           ,x"c060"
           ,x"600e"
           ,x"0281"
           ,x"6072"
           ,x"1602"
           ,x"0460"
           ,x"6072"
           ,x"0420"
           ,x"000c"
           ,x"18ef"
           ,x"0204"
           ,x"0003"
           ,x"04c0"
           ,x"d800"
           ,x"9c02"
           ,x"06c0"
           ,x"d800"
           ,x"9c02"
           ,x"06c0"
           ,x"c800"
           ,x"8322"
           ,x"0420"
           ,x"0010"
           ,x"04c1"
           ,x"0202"
           ,x"1800"
           ,x"04c3"
           ,x"d0e0"
           ,x"9800"
           ,x"0b11"
           ,x"a043"
           ,x"0602"
           ,x"16f9"
           ,x"c801"
           ,x"8322"
           ,x"0420"
           ,x"0010"
           ,x"04c1"
           ,x"d060"
           ,x"9802"
           ,x"d0a0"
           ,x"9802"
           ,x"0982"
           ,x"e042"
           ,x"c801"
           ,x"8322"
           ,x"0420"
           ,x"0010"
           ,x"0420"
           ,x"000c"
           ,x"0524"
           ,x"0220"
           ,x"2000"
           ,x"0280"
           ,x"6000"
           ,x"16d5"
           ,x"0604"
           ,x"16d2"
           ,x"0420"
           ,x"001c"
           ,x"102c"
           ,x"0202"
           ,x"04fc"
           ,x"0201"
           ,x"0020"
           ,x"0203"
           ,x"4300"
           ,x"06c3"
           ,x"d803"
           ,x"8c02"
           ,x"06c3"
           ,x"d803"
           ,x"8c02"
           ,x"d832"
           ,x"8c00"
           ,x"0601"
           ,x"16fc"
           ,x"0203"
           ,x"4000"
           ,x"06c3"
           ,x"d803"
           ,x"8c02"
           ,x"06c3"
           ,x"d803"
           ,x"8c02"
           ,x"0205"
           ,x"0080"
           ,x"0200"
           ,x"2021"
           ,x"d800"
           ,x"8c00"
           ,x"06c0"
           ,x"d800"
           ,x"8c00"
           ,x"06c0"
           ,x"0200"
           ,x"3031"
           ,x"d800"
           ,x"8c00"
           ,x"06c0"
           ,x"d800"
           ,x"8c00"
           ,x"06c0"
           ,x"0605"
           ,x"16ee"
           ,x"0201"
           ,x"b000"
           ,x"0200"
           ,x"0100"
           ,x"0203"
           ,x"0014"
           ,x"d440"
           ,x"0a10"
           ,x"1602"
           ,x"0200"
           ,x"0100"
           ,x"04c2"
           ,x"0602"
           ,x"16fe"
           ,x"0603"
           ,x"16f6"
           ,x"0200"
           ,x"0000"
           ,x"06a0"
           ,x"038a"
           ,x"0201"
           ,x"0dc0"
           ,x"0202"
           ,x"0b10"
           ,x"d831"
           ,x"8c00"
           ,x"d831"
           ,x"8c00"
           ,x"0642"
           ,x"16fa"
           ,x"0201"
           ,x"000a"
           ,x"0602"
           ,x"16fe"
           ,x"0601"
           ,x"16fc"
           ,x"0204"
           ,x"10a0"
           ,x"0205"
           ,x"0000"
           ,x"0206"
           ,x"0000"
           ,x"0208"
           ,x"0020"
           ,x"c081"
           ,x"0209"
           ,x"2710"
           ,x"0201"
           ,x"0dc0"
           ,x"04c0"
           ,x"06a0"
           ,x"038a"
           ,x"c1c6"
           ,x"a1c5"
           ,x"0247"
           ,x"001f"
           ,x"a1c1"
           ,x"d817"
           ,x"8c00"
           ,x"0586"
           ,x"8206"
           ,x"16f6"
           ,x"04c6"
           ,x"0221"
           ,x"0020"
           ,x"8101"
           ,x"16f1"
           ,x"0585"
           ,x"0245"
           ,x"001f"
           ,x"0289"
           ,x"0000"
           ,x"13e6"
           ,x"c1c9"
           ,x"0607"
           ,x"16fe"
           ,x"0229"
           ,x"fff6"
           ,x"0200"
           ,x"02e0"
           ,x"c800"
           ,x"8320"
           ,x"0420"
           ,x"000c"
           ,x"18d0"
           ,x"c809"
           ,x"8322"
           ,x"0420"
           ,x"0010"
           ,x"0420"
           ,x"000c"
           ,x"18ec"
           ,x"0221"
           ,x"0020"
           ,x"10d0"
           ,x"10a0"
           ,x"0240"
           ,x"3fff"
           ,x"06c0"
           ,x"d800"
           ,x"8c02"
           ,x"06c0"
           ,x"0260"
           ,x"4000"
           ,x"d800"
           ,x"8c02"
           ,x"045b"
           ,x"c28b"
           ,x"0206"
           ,x"0020"
           ,x"04c0"
           ,x"0207"
           ,x"0017"
           ,x"06c6"
           ,x"d806"
           ,x"8c02"
           ,x"06c6"
           ,x"d806"
           ,x"8c02"
           ,x"0202"
           ,x"0020"
           ,x"0205"
           ,x"a040"
           ,x"0201"
           ,x"8800"
           ,x"dd51"
           ,x"dd51"
           ,x"0642"
           ,x"16fc"
           ,x"06a0"
           ,x"038a"
           ,x"0202"
           ,x"0020"
           ,x"0205"
           ,x"a040"
           ,x"0201"
           ,x"8c00"
           ,x"d475"
           ,x"d475"
           ,x"0642"
           ,x"16fc"
           ,x"0220"
           ,x"0020"
           ,x"0226"
           ,x"0020"
           ,x"0607"
           ,x"16de"
           ,x"045a"
           ,x"c28b"
           ,x"0200"
           ,x"06b4"
           ,x"0207"
           ,x"0528"
           ,x"a1c0"
           ,x"0200"
           ,x"0900"
           ,x"06a0"
           ,x"038a"
           ,x"0200"
           ,x"003e"
           ,x"04c2"
           ,x"0201"
           ,x"0007"
           ,x"d837"
           ,x"8c00"
           ,x"0601"
           ,x"16fc"
           ,x"d802"
           ,x"8c00"
           ,x"0600"
           ,x"16f6"
           ,x"045a"
           ,x"0203"
           ,x"0004"
           ,x"c28b"
           ,x"c081"
           ,x"06a0"
           ,x"043e"
           ,x"0a42"
           ,x"c042"
           ,x"0603"
           ,x"16fa"
           ,x"045a"
           ,x"0203"
           ,x"0002"
           ,x"10f4"
           ,x"0941"
           ,x"0241"
           ,x"0f00"
           ,x"0221"
           ,x"3000"
           ,x"0281"
           ,x"3a00"
           ,x"1a02"
           ,x"0221"
           ,x"0700"
           ,x"d801"
           ,x"8c00"
           ,x"045b"
           ,x"0300"
           ,x"0000"
           ,x"06a0"
           ,x"038a"
           ,x"06a0"
           ,x"0422"
           ,x"0220"
           ,x"0004"
           ,x"0380"
           ,x"0300"
           ,x"0000"
           ,x"c07e"
           ,x"06a0"
           ,x"038a"
           ,x"d0b1"
           ,x"1311"
           ,x"0282"
           ,x"0d00"
           ,x"13fb"
           ,x"0282"
           ,x"0a00"
           ,x"1607"
           ,x"0220"
           ,x"0020"
           ,x"0240"
           ,x"ffe0"
           ,x"06a0"
           ,x"038a"
           ,x"10f1"
           ,x"0580"
           ,x"d802"
           ,x"8c00"
           ,x"10ed"
           ,x"0380"
           ,x"0300"
           ,x"0000"
           ,x"06a0"
           ,x"038a"
           ,x"0580"
           ,x"d801"
           ,x"8c00"
           ,x"0380"
           ,x"0300"
           ,x"0000"
           ,x"04c0"
           ,x"0201"
           ,x"2000"
           ,x"0202"
           ,x"0300"
           ,x"d820"
           ,x"8321"
           ,x"8c02"
           ,x"0260"
           ,x"4000"
           ,x"d800"
           ,x"8c02"
           ,x"d801"
           ,x"8c00"
           ,x"0602"
           ,x"16fc"
           ,x"0200"
           ,x"0001"
           ,x"06a0"
           ,x"038a"
           ,x"0380"
           ,x"04c0"
           ,x"0201"
           ,x"000a"
           ,x"0600"
           ,x"16fe"
           ,x"0601"
           ,x"16fc"
           ,x"06a0"
           ,x"03a0"
           ,x"04c0"
           ,x"0201"
           ,x"000a"
           ,x"0600"
           ,x"16fe"
           ,x"0601"
           ,x"16fc"
           ,x"0380"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0018"
           ,x"2442"
           ,x"427e"
           ,x"4242"
           ,x"8080"
           ,x"8080"
           ,x"8080"
           ,x"8080"
           ,x"0103"
           ,x"0101"
           ,x"0101"
           ,x"0101"
           ,x"00e0"
           ,x"000e"
           ,x"0106"
           ,x"00f7"
           ,x"0d0a"
           ,x"0000"
           ,x"aa02"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"1310"
           ,x"1320"
           ,x"0000"
           ,x"0000"
           ,x"43dc"
           ,x"443c"
           ,x"49a9"
           ,x"4396"
           ,x"439e"
           ,x"4446"
           ,x"4449"
           ,x"444c"
           ,x"4052"
           ,x"51fe"
           ,x"4c82"
           ,x"4d59"
           ,x"4db4"
           ,x"4e64"
           ,x"4ef9"
           ,x"4f01"
           ,x"4f5f"
           ,x"4f80"
           ,x"43ce"
           ,x"43d6"
           ,x"054d"
           ,x"1252"
           ,x"5e44"
           ,x"1705"
           ,x"2844"
           ,x"0537"
           ,x"b460"
           ,x"0d00"
           ,x"1100"
           ,x"43c2"
           ,x"04b4"
           ,x"06b4"
           ,x"0874"
           ,x"8780"
           ,x"cebe"
           ,x"8f11"
           ,x"0070"
           ,x"be81"
           ,x"009f"
           ,x"be81"
           ,x"00bf"
           ,x"be81"
           ,x"00df"
           ,x"be81"
           ,x"00ff"
           ,x"bf72"
           ,x"ff7e"
           ,x"3900"
           ,x"0800"
           ,x"0451"
           ,x"8600"
           ,x"3500"
           ,x"7101"
           ,x"0035"
           ,x"003e"
           ,x"8082"
           ,x"0035"
           ,x"000b"
           ,x"7400"
           ,x"3500"
           ,x"0880"
           ,x"c200"
           ,x"bf03"
           ,x"0308"
           ,x"f602"
           ,x"03bf"
           ,x"0310"
           ,x"01f6"
           ,x"0203"
           ,x"be03"
           ,x"18f6"
           ,x"0203"
           ,x"8400"
           ,x"be03"
           ,x"02f6"
           ,x"0203"
           ,x"be03"
           ,x"01f6"
           ,x"0203"
           ,x"bf03"
           ,x"1602"
           ,x"f602"
           ,x"0306"
           ,x"03ce"
           ,x"86a0"
           ,x"00be"
           ,x"7010"
           ,x"beb0"
           ,x"70a0"
           ,x"8ea0"
           ,x"0040"
           ,x"dc39"
           ,x"0001"
           ,x"0104"
           ,x"4f86"
           ,x"b070"
           ,x"a070"
           ,x"70d6"
           ,x"7040"
           ,x"40be"
           ,x"be80"
           ,x"fd08"
           ,x"9370"
           ,x"3900"
           ,x"0101"
           ,x"0244"
           ,x"86a0"
           ,x"0035"
           ,x"0fff"
           ,x"a001"
           ,x"a000"
           ,x"3100"
           ,x"20a3"
           ,x"8004"
           ,x"5931"
           ,x"0200"
           ,x"a900"
           ,x"04b4"
           ,x"3100"
           ,x"50a8"
           ,x"0809"
           ,x"5007"
           ,x"20be"
           ,x"7e05"
           ,x"bc74"
           ,x"7e03"
           ,x"927e"
           ,x"4108"
           ,x"877e"
           ,x"be75"
           ,x"6008"
           ,x"c1e0"
           ,x"75fb"
           ,x"0117"
           ,x"b09d"
           ,x"c1e0"
           ,x"75fb"
           ,x"011f"
           ,x"fba6"
           ,x"7e12"
           ,x"a275"
           ,x"08d6"
           ,x"75e0"
           ,x"4115"
           ,x"d67e"
           ,x"0341"
           ,x"1287"
           ,x"7e08"
           ,x"a48e"
           ,x"0201"
           ,x"0203"
           ,x"9c02"
           ,x"0405"
           ,x"069c"
           ,x"0207"
           ,x"0809"
           ,x"a78f"
           ,x"1b52"
           ,x"4541"
           ,x"4459"
           ,x"2d50"
           ,x"5245"
           ,x"5353"
           ,x"2041"
           ,x"4e59"
           ,x"204b"
           ,x"4559"
           ,x"2054"
           ,x"4f20"
           ,x"4245"
           ,x"4749"
           ,x"4efb"
           ,x"3100"
           ,x"11a1"
           ,x"2804"
           ,x"9631"
           ,x"0018"
           ,x"a2c4"
           ,x"048f"
           ,x"3100"
           ,x"0da1"
           ,x"6a04"
           ,x"a7be"
           ,x"4310"
           ,x"0603"
           ,x"7c87"
           ,x"80d0"
           ,x"8655"
           ,x"be6d"
           ,x"040f"
           ,x"1961"
           ,x"8bbf"
           ,x"7200"
           ,x"80bf"
           ,x"9072"
           ,x"01a2"
           ,x"0f1a"
           ,x"bd90"
           ,x"7390"
           ,x"7296"
           ,x"7200"
           ,x"8f80"
           ,x"d041"
           ,x"8f39"
           ,x"0001"
           ,x"0104"
           ,x"5086"
           ,x"7402"
           ,x"ff03"
           ,x"41af"
           ,x"0603"
           ,x"ce07"
           ,x"20be"
           ,x"72fe"
           ,x"be6d"
           ,x"0686"
           ,x"6c86"
           ,x"80fb"
           ,x"3100"
           ,x"1ea4"
           ,x"0060"
           ,x"00be"
           ,x"80fb"
           ,x"0431"
           ,x"001e"
           ,x"a420"
           ,x"6000"
           ,x"8658"
           ,x"8659"
           ,x"0501"
           ,x"df90"
           ,x"59ce"
           ,x"591d"
           ,x"61f0"
           ,x"d4e4"
           ,x"0058"
           ,x"e420"
           ,x"5841"
           ,x"f205"
           ,x"01dd"
           ,x"4200"
           ,x"9472"
           ,x"8790"
           ,x"7294"
           ,x"72bf"
           ,x"9072"
           ,x"12a5"
           ,x"906c"
           ,x"d68f"
           ,x"dd00"
           ,x"aa42"
           ,x"27bd"
           ,x"588f"
           ,x"dd06"
           ,x"8f58"
           ,x"6227"
           ,x"9472"
           ,x"bf90"
           ,x"72ff"
           ,x"ff94"
           ,x"72bd"
           ,x"9072"
           ,x"5890"
           ,x"6cbd"
           ,x"58cf"
           ,x"7d00"
           ,x"5842"
           ,x"0c94"
           ,x"7287"
           ,x"9072"
           ,x"0f1a"
           ,x"6227"
           ,x"9672"
           ,x"d702"
           ,x"12a5"
           ,x"4243"
           ,x"3100"
           ,x"0159"
           ,x"6000"
           ,x"d659"
           ,x"aa41"
           ,x"b939"
           ,x"0001"
           ,x"0104"
           ,x"5108"
           ,x"a081"
           ,x"0201"
           ,x"0203"
           ,x"9c02"
           ,x"0405"
           ,x"069c"
           ,x"0207"
           ,x"0809"
           ,x"a09e"
           ,x"0450"
           ,x"5245"
           ,x"5353"
           ,x"fb31"
           ,x"0011"
           ,x"a028"
           ,x"0496"
           ,x"3100"
           ,x"0da0"
           ,x"6804"
           ,x"a7bf"
           ,x"5200"
           ,x"e4be"
           ,x"5830"
           ,x"8e6c"
           ,x"4293"
           ,x"08ff"
           ,x"020f"
           ,x"494e"
           ,x"5345"
           ,x"5254"
           ,x"2043"
           ,x"4152"
           ,x"5452"
           ,x"4944"
           ,x"4745"
           ,x"fb42"
           ,x"ef90"
           ,x"58bc"
           ,x"b052"
           ,x"5895"
           ,x"5231"
           ,x"0003"
           ,x"b052"
           ,x"094d"
           ,x"a352"
           ,x"0004"
           ,x"bd6a"
           ,x"9072"
           ,x"9672"
           ,x"bd5c"
           ,x"9072"
           ,x"9672"
           ,x"a36a"
           ,x"0004"
           ,x"865e"
           ,x"8e5c"
           ,x"62d0"
           ,x"3500"
           ,x"015f"
           ,x"cf7d"
           ,x"006a"
           ,x"916a"
           ,x"345e"
           ,x"b052"
           ,x"cf7d"
           ,x"006a"
           ,x"42e0"
           ,x"3300"
           ,x"015f"
           ,x"0000"
           ,x"6a91"
           ,x"6a32"
           ,x"5eb0"
           ,x"5200"
           ,x"006a"
           ,x"a352"
           ,x"003a"
           ,x"d272"
           ,x"0062"
           ,x"93be"
           ,x"4313"
           ,x"0603"
           ,x"7c39"
           ,x"0001"
           ,x"0104"
           ,x"5086"
           ,x"7402"
           ,x"ff03"
           ,x"42f7"
           ,x"a675"
           ,x"31c8"
           ,x"756c"
           ,x"430a"
           ,x"0603"
           ,x"d605"
           ,x"02f7"
           ,x"0603"
           ,x"cea4"
           ,x"6c75"
           ,x"926c"
           ,x"e26c"
           ,x"02bc"
           ,x"7890"
           ,x"6c94"
           ,x"6cbd"
           ,x"5c90"
           ,x"6c95"
           ,x"5cbf"
           ,x"729e"
           ,x"808e"
           ,x"7863"
           ,x"32bd"
           ,x"8080"
           ,x"cf7d"
           ,x"005c"
           ,x"433a"
           ,x"3300"
           ,x"0280"
           ,x"8000"
           ,x"005c"
           ,x"0720"
           ,x"8f80"
           ,x"ce43"
           ,x"3ccf"
           ,x"7010"
           ,x"0043"
           ,x"56bd"
           ,x"0070"
           ,x"a700"
           ,x"0fff"
           ,x"3400"
           ,x"af10"
           ,x"00af"
           ,x"0fff"
           ,x"8600"
           ,x"3500"
           ,x"6f01"
           ,x"0035"
           ,x"003c"
           ,x"8084"
           ,x"0086"
           ,x"7435"
           ,x"001f"
           ,x"a381"
           ,x"a380"
           ,x"8780"
           ,x"828e"
           ,x"7863"
           ,x"7b96"
           ,x"73bd"
           ,x"0080"
           ,x"800f"
           ,x"f000"
           ,x"be42"
           ,x"6031"
           ,x"0002"
           ,x"2860"
           ,x"00d6"
           ,x"28aa"
           ,x"4395"
           ,x"d229"
           ,x"0063"
           ,x"9594"
           ,x"73bd"
           ,x"9073"
           ,x"4200"
           ,x"3102"
           ,x"00b0"
           ,x"4a04"
           ,x"b400"
           ,x"bf80"
           ,x"d006"
           ,x"b4be"
           ,x"80d2"
           ,x"4086"
           ,x"b04a"
           ,x"3300"
           ,x"07e0"
           ,x"014a"
           ,x"0000"
           ,x"d0a3"
           ,x"4a00"
           ,x"08a3"
           ,x"80d0"
           ,x"0007"
           ,x"9280"
           ,x"d243"
           ,x"a700"
           ,x"bf80"
           ,x"d008"
           ,x"74be"
           ,x"80d2"
           ,x"1f05"
           ,x"03a7"
           ,x"bf58"
           ,x"0479"
           ,x"f658"
           ,x"0000"
           ,x"bf58"
           ,x"0484"
           ,x"43d2"
           ,x"886d"
           ,x"8654"
           ,x"bc55"
           ,x"b056"
           ,x"8658"
           ,x"bd52"
           ,x"5691"
           ,x"52d4"
           ,x"5855"
           ,x"63fa"
           ,x"d6b0"
           ,x"522e"
           ,x"63fa"
           ,x"9058"
           ,x"43e9"
           ,x"8e58"
           ,x"6438"
           ,x"bc55"
           ,x"58d2"
           ,x"5508"
           ,x"6438"
           ,x"8654"
           ,x"8780"
           ,x"d091"
           ,x"5634"
           ,x"544a"
           ,x"b056"
           ,x"a156"
           ,x"540f"
           ,x"1994"
           ,x"73bd"
           ,x"9073"
           ,x"80fa"
           ,x"0f1a"
           ,x"442c"
           ,x"9473"
           ,x"bd90"
           ,x"7390"
           ,x"7296"
           ,x"7200"
           ,x"8f80"
           ,x"d044"
           ,x"1ebd"
           ,x"80fa"
           ,x"9073"
           ,x"9673"
           ,x"d400"
           ,x"0001"
           ,x"9673"
           ,x"bd80"
           ,x"fa90"
           ,x"7396"
           ,x"7300"
           ,x"0528"
           ,x"4c05"
           ,x"284e"
           ,x"0520"
           ,x"1080"
           ,x"6000"
           ,x"20f0"
           ,x"0ef9"
           ,x"86f8"
           ,x"f717"
           ,x"1717"
           ,x"1717"
           ,x"1717"
           ,x"1717"
           ,x"1717"
           ,x"1706"
           ,x"0301"
           ,x"0b0c"
           ,x"0d0f"
           ,x"0402"
           ,x"0d08"
           ,x"0e05"
           ,x"090a"
           ,x"0627"
           ,x"2722"
           ,x"2206"
           ,x"bfdf"
           ,x"ff80"
           ,x"0592"
           ,x"0a01"
           ,x"9f00"
           ,x"06bf"
           ,x"dfff"
           ,x"8020"
           ,x"900a"
           ,x"019f"
           ,x"000a"
           ,x"3139"
           ,x"3831"
           ,x"2020"
           ,x"5445"
           ,x"5841"
           ,x"5320"
           ,x"494e"
           ,x"5354"
           ,x"5255"
           ,x"4d45"
           ,x"4e54"
           ,x"5348"
           ,x"4f4d"
           ,x"4520"
           ,x"434f"
           ,x"4d50"
           ,x"5554"
           ,x"4552"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"0020"
           ,x"4848"
           ,x"4800"
           ,x"0000"
           ,x"0000"
           ,x"0048"
           ,x"fc48"
           ,x"48fc"
           ,x"4800"
           ,x"103c"
           ,x"5038"
           ,x"1478"
           ,x"1000"
           ,x"c0c4"
           ,x"0810"
           ,x"2040"
           ,x"8c0c"
           ,x"6090"
           ,x"9060"
           ,x"6094"
           ,x"8874"
           ,x"0810"
           ,x"2000"
           ,x"0000"
           ,x"0000"
           ,x"0810"
           ,x"2020"
           ,x"2020"
           ,x"1008"
           ,x"4020"
           ,x"1010"
           ,x"1010"
           ,x"2040"
           ,x"0000"
           ,x"4830"
           ,x"cc30"
           ,x"4800"
           ,x"0000"
           ,x"1010"
           ,x"7c10"
           ,x"1000"
           ,x"0000"
           ,x"0000"
           ,x"0030"
           ,x"1020"
           ,x"0000"
           ,x"0000"
           ,x"7c00"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"3030"
           ,x"0004"
           ,x"0810"
           ,x"2040"
           ,x"8000"
           ,x"3844"
           ,x"4444"
           ,x"4444"
           ,x"4438"
           ,x"1030"
           ,x"5010"
           ,x"1010"
           ,x"107c"
           ,x"7884"
           ,x"0408"
           ,x"1020"
           ,x"40fc"
           ,x"7884"
           ,x"0438"
           ,x"0404"
           ,x"8478"
           ,x"0c14"
           ,x"2444"
           ,x"84fc"
           ,x"0404"
           ,x"f880"
           ,x"80f8"
           ,x"0404"
           ,x"8478"
           ,x"7880"
           ,x"80f8"
           ,x"8484"
           ,x"8478"
           ,x"fc04"
           ,x"0408"
           ,x"1020"
           ,x"4040"
           ,x"7884"
           ,x"8478"
           ,x"8484"
           ,x"8478"
           ,x"7884"
           ,x"8484"
           ,x"7c04"
           ,x"0478"
           ,x"0030"
           ,x"3000"
           ,x"0030"
           ,x"3000"
           ,x"0030"
           ,x"3000"
           ,x"0030"
           ,x"1020"
           ,x"0008"
           ,x"1020"
           ,x"4020"
           ,x"1008"
           ,x"0000"
           ,x"007c"
           ,x"007c"
           ,x"0000"
           ,x"0040"
           ,x"2010"
           ,x"0810"
           ,x"2040"
           ,x"3844"
           ,x"0408"
           ,x"1010"
           ,x"0010"
           ,x"0078"
           ,x"849c"
           ,x"a498"
           ,x"807c"
           ,x"7884"
           ,x"8484"
           ,x"fc84"
           ,x"8484"
           ,x"f844"
           ,x"4478"
           ,x"4444"
           ,x"44f8"
           ,x"7884"
           ,x"8080"
           ,x"8080"
           ,x"8478"
           ,x"f844"
           ,x"4444"
           ,x"4444"
           ,x"44f8"
           ,x"fc80"
           ,x"80f0"
           ,x"8080"
           ,x"80fc"
           ,x"fc80"
           ,x"80f0"
           ,x"8080"
           ,x"8080"
           ,x"7884"
           ,x"8080"
           ,x"9c84"
           ,x"8478"
           ,x"8484"
           ,x"84fc"
           ,x"8484"
           ,x"8484"
           ,x"7c10"
           ,x"1010"
           ,x"1010"
           ,x"107c"
           ,x"0404"
           ,x"0404"
           ,x"0484"
           ,x"8478"
           ,x"8890"
           ,x"a0c0"
           ,x"a090"
           ,x"8884"
           ,x"4040"
           ,x"4040"
           ,x"4040"
           ,x"407c"
           ,x"84cc"
           ,x"b484"
           ,x"8484"
           ,x"8484"
           ,x"84c4"
           ,x"a494"
           ,x"8c84"
           ,x"8484"
           ,x"fc84"
           ,x"8484"
           ,x"8484"
           ,x"84fc"
           ,x"f884"
           ,x"8484"
           ,x"f880"
           ,x"8080"
           ,x"7884"
           ,x"8484"
           ,x"8494"
           ,x"8874"
           ,x"f884"
           ,x"8484"
           ,x"f890"
           ,x"8884"
           ,x"7884"
           ,x"8078"
           ,x"0404"
           ,x"8478"
           ,x"7c10"
           ,x"1010"
           ,x"1010"
           ,x"1010"
           ,x"8484"
           ,x"8484"
           ,x"8484"
           ,x"8478"
           ,x"4444"
           ,x"4444"
           ,x"2828"
           ,x"1010"
           ,x"8484"
           ,x"8484"
           ,x"84b4"
           ,x"cc84"
           ,x"8484"
           ,x"4830"
           ,x"3048"
           ,x"8484"
           ,x"4444"
           ,x"4428"
           ,x"1010"
           ,x"1010"
           ,x"fc04"
           ,x"0810"
           ,x"2040"
           ,x"80fc"
           ,x"3820"
           ,x"2020"
           ,x"2020"
           ,x"2038"
           ,x"0080"
           ,x"4020"
           ,x"1008"
           ,x"0400"
           ,x"7010"
           ,x"1010"
           ,x"1010"
           ,x"1070"
           ,x"1028"
           ,x"4482"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"00fc"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0010"
           ,x"1010"
           ,x"1010"
           ,x"0010"
           ,x"2828"
           ,x"2800"
           ,x"0000"
           ,x"0028"
           ,x"287c"
           ,x"287c"
           ,x"2828"
           ,x"3854"
           ,x"5038"
           ,x"1454"
           ,x"3860"
           ,x"6408"
           ,x"1020"
           ,x"4c0c"
           ,x"2050"
           ,x"5020"
           ,x"5448"
           ,x"3408"
           ,x"0810"
           ,x"0000"
           ,x"0000"
           ,x"0810"
           ,x"2020"
           ,x"2010"
           ,x"0820"
           ,x"1008"
           ,x"0808"
           ,x"1020"
           ,x"0028"
           ,x"107c"
           ,x"1028"
           ,x"0000"
           ,x"1010"
           ,x"7c10"
           ,x"1000"
           ,x"0000"
           ,x"0000"
           ,x"3010"
           ,x"2000"
           ,x"0000"
           ,x"7c00"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0030"
           ,x"3000"
           ,x"0408"
           ,x"1020"
           ,x"4000"
           ,x"3844"
           ,x"4444"
           ,x"4444"
           ,x"3810"
           ,x"3010"
           ,x"1010"
           ,x"1038"
           ,x"3844"
           ,x"0408"
           ,x"1020"
           ,x"7c38"
           ,x"4404"
           ,x"1804"
           ,x"4438"
           ,x"0818"
           ,x"2848"
           ,x"7c08"
           ,x"087c"
           ,x"4078"
           ,x"0404"
           ,x"4438"
           ,x"1820"
           ,x"4078"
           ,x"4444"
           ,x"387c"
           ,x"0408"
           ,x"1020"
           ,x"2020"
           ,x"3844"
           ,x"4438"
           ,x"4444"
           ,x"3838"
           ,x"4444"
           ,x"3c04"
           ,x"0830"
           ,x"0030"
           ,x"3000"
           ,x"3030"
           ,x"0000"
           ,x"3030"
           ,x"0030"
           ,x"1020"
           ,x"0810"
           ,x"2040"
           ,x"2010"
           ,x"0800"
           ,x"007c"
           ,x"007c"
           ,x"0000"
           ,x"2010"
           ,x"0804"
           ,x"0810"
           ,x"2038"
           ,x"4404"
           ,x"0810"
           ,x"0010"
           ,x"3844"
           ,x"5c54"
           ,x"5c40"
           ,x"3838"
           ,x"4444"
           ,x"7c44"
           ,x"4444"
           ,x"7824"
           ,x"2438"
           ,x"2424"
           ,x"7838"
           ,x"4440"
           ,x"4040"
           ,x"4438"
           ,x"7824"
           ,x"2424"
           ,x"2424"
           ,x"787c"
           ,x"4040"
           ,x"7840"
           ,x"407c"
           ,x"7c40"
           ,x"4078"
           ,x"4040"
           ,x"403c"
           ,x"4040"
           ,x"5c44"
           ,x"4438"
           ,x"4444"
           ,x"447c"
           ,x"4444"
           ,x"4438"
           ,x"1010"
           ,x"1010"
           ,x"1038"
           ,x"0404"
           ,x"0404"
           ,x"0444"
           ,x"3844"
           ,x"4850"
           ,x"6050"
           ,x"4844"
           ,x"4040"
           ,x"4040"
           ,x"4040"
           ,x"7c44"
           ,x"6c54"
           ,x"5444"
           ,x"4444"
           ,x"4464"
           ,x"6454"
           ,x"4c4c"
           ,x"447c"
           ,x"4444"
           ,x"4444"
           ,x"447c"
           ,x"7844"
           ,x"4478"
           ,x"4040"
           ,x"4038"
           ,x"4444"
           ,x"4454"
           ,x"4834"
           ,x"7844"
           ,x"4478"
           ,x"5048"
           ,x"4438"
           ,x"4440"
           ,x"3804"
           ,x"4438"
           ,x"7c10"
           ,x"1010"
           ,x"1010"
           ,x"1044"
           ,x"4444"
           ,x"4444"
           ,x"4438"
           ,x"4444"
           ,x"4428"
           ,x"2810"
           ,x"1044"
           ,x"4444"
           ,x"5454"
           ,x"5428"
           ,x"4444"
           ,x"2810"
           ,x"2844"
           ,x"4444"
           ,x"4428"
           ,x"1010"
           ,x"1010"
           ,x"7c04"
           ,x"0810"
           ,x"2040"
           ,x"7c38"
           ,x"2020"
           ,x"2020"
           ,x"2038"
           ,x"0040"
           ,x"2010"
           ,x"0804"
           ,x"0038"
           ,x"0808"
           ,x"0808"
           ,x"0838"
           ,x"0010"
           ,x"2844"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"007c"
           ,x"0020"
           ,x"1008"
           ,x"0000"
           ,x"0000"
           ,x"0038"
           ,x"447c"
           ,x"4444"
           ,x"0000"
           ,x"7824"
           ,x"3824"
           ,x"7800"
           ,x"003c"
           ,x"4040"
           ,x"403c"
           ,x"0000"
           ,x"7824"
           ,x"2424"
           ,x"7800"
           ,x"6060"
           ,x"6868"
           ,x"7070"
           ,x"7878"
           ,x"8080"
           ,x"8888"
           ,x"9090"
           ,x"9898"
           ,x"a0a0"
           ,x"a8a8"
           ,x"b0b0"
           ,x"b8b8"
           ,x"c0c0"
           ,x"c8c8"
           ,x"d0d0"
           ,x"d8d8"
           ,x"6060"
           ,x"6868"
           ,x"7070"
           ,x"7878"
           ,x"8080"
           ,x"8888"
           ,x"9090"
           ,x"9898"
           ,x"a0a0"
           ,x"a8a8"
           ,x"b0b0"
           ,x"b8b8"
           ,x"c0c0"
           ,x"c8c8"
           ,x"d0d0"
           ,x"d8d8"
           ,x"6060"
           ,x"6868"
           ,x"7070"
           ,x"7878"
           ,x"8080"
           ,x"8888"
           ,x"9090"
           ,x"9898"
           ,x"a0a0"
           ,x"a8a8"
           ,x"b0b0"
           ,x"b8b8"
           ,x"c0c0"
           ,x"c8c8"
           ,x"d0d0"
           ,x"d8d8"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2001"
           ,x"0203"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2004"
           ,x"0506"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2007"
           ,x"0809"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"5445"
           ,x"5841"
           ,x"5320"
           ,x"494e"
           ,x"5354"
           ,x"5255"
           ,x"4d45"
           ,x"4e54"
           ,x"5320"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"484f"
           ,x"4d45"
           ,x"2043"
           ,x"4f4d"
           ,x"5055"
           ,x"5445"
           ,x"5220"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"5245"
           ,x"4144"
           ,x"592d"
           ,x"5052"
           ,x"4553"
           ,x"5320"
           ,x"414e"
           ,x"5920"
           ,x"4b45"
           ,x"5920"
           ,x"544f"
           ,x"2042"
           ,x"4547"
           ,x"494e"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"6060"
           ,x"6868"
           ,x"7070"
           ,x"7878"
           ,x"8080"
           ,x"8888"
           ,x"9090"
           ,x"9898"
           ,x"a0a0"
           ,x"a8a8"
           ,x"b0b0"
           ,x"b8b8"
           ,x"c0c0"
           ,x"c8c8"
           ,x"d0d0"
           ,x"d8d8"
           ,x"6060"
           ,x"6868"
           ,x"7070"
           ,x"7878"
           ,x"8080"
           ,x"8888"
           ,x"9090"
           ,x"9898"
           ,x"a0a0"
           ,x"a8a8"
           ,x"b0b0"
           ,x"b8b8"
           ,x"c0c0"
           ,x"c8c8"
           ,x"d0d0"
           ,x"d8d8"
           ,x"6060"
           ,x"6868"
           ,x"7070"
           ,x"7878"
           ,x"8080"
           ,x"8888"
           ,x"9090"
           ,x"9898"
           ,x"a0a0"
           ,x"a8a8"
           ,x"b0b0"
           ,x"b8b8"
           ,x"c0c0"
           ,x"c8c8"
           ,x"d0d0"
           ,x"d8d8"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"0a31"
           ,x"3938"
           ,x"3120"
           ,x"2054"
           ,x"4558"
           ,x"4153"
           ,x"2049"
           ,x"4e53"
           ,x"5452"
           ,x"554d"
           ,x"454e"
           ,x"5453"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"1717"
           ,x"1717"
           ,x"1717"
           ,x"1717"
           ,x"1717"
           ,x"1717"
           ,x"0603"
           ,x"010b"
           ,x"0c0d"
           ,x"0f04"
           ,x"020d"
           ,x"080e"
           ,x"0509"
           ,x"0a06"
           ,x"2727"
           ,x"2222"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0103"
           ,x"0303"
           ,x"0303"
           ,x"0303"
           ,x"fc04"
           ,x"0505"
           ,x"0406"
           ,x"020c"
           ,x"0080"
           ,x"4040"
           ,x"8000"
           ,x"0c12"
           ,x"ff80"
           ,x"c040"
           ,x"6038"
           ,x"1c0e"
           ,x"1921"
           ,x"213d"
           ,x"0505"
           ,x"05c4"
           ,x"ba8a"
           ,x"8aba"
           ,x"a1a1"
           ,x"a122"
           ,x"0301"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"e231"
           ,x"1018"
           ,x"0c07"
           ,x"0300"
           ,x"4c90"
           ,x"2040"
           ,x"4020"
           ,x"e000"
           ,x"3c42"
           ,x"99a1"
           ,x"a199"
           ,x"423c"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"2020"
           ,x"2020"
           ,x"2020"
           ,x"0020"
           ,x"4848"
           ,x"4800"
           ,x"0000"
           ,x"0000"
           ,x"0048"
           ,x"fc48"
           ,x"48fc"
           ,x"4800"
           ,x"103c"
           ,x"5038"
           ,x"1478"
           ,x"1000"
           ,x"c0c4"
           ,x"0810"
           ,x"2040"
           ,x"8c0c"
           ,x"6090"
           ,x"9060"
           ,x"6094"
           ,x"8874"
           ,x"0810"
           ,x"2000"
           ,x"0000"
           ,x"0000"
           ,x"0810"
           ,x"2020"
           ,x"2020"
           ,x"1008"
           ,x"4020"
           ,x"1010"
           ,x"1010"
           ,x"2040"
           ,x"0000"
           ,x"4830"
           ,x"cc30"
           ,x"4800"
           ,x"0000"
           ,x"1010"
           ,x"7c10"
           ,x"1000"
           ,x"0000"
           ,x"0000"
           ,x"0030"
           ,x"1020"
           ,x"0000"
           ,x"0000"
           ,x"7c00"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"3030"
           ,x"0004"
           ,x"0810"
           ,x"2040"
           ,x"8000"
           ,x"3844"
           ,x"4444"
           ,x"4444"
           ,x"4438"
           ,x"1030"
           ,x"5010"
           ,x"1010"
           ,x"107c"
           ,x"7884"
           ,x"0408"
           ,x"1020"
           ,x"40fc"
           ,x"7884"
           ,x"0438"
           ,x"0404"
           ,x"8478"
           ,x"0c14"
           ,x"2444"
           ,x"84fc"
           ,x"0404"
           ,x"f880"
           ,x"80f8"
           ,x"0404"
           ,x"8478"
           ,x"7880"
           ,x"80f8"
           ,x"8484"
           ,x"8478"
           ,x"fc04"
           ,x"0408"
           ,x"1020"
           ,x"4040"
           ,x"7884"
           ,x"8478"
           ,x"8484"
           ,x"8478"
           ,x"7884"
           ,x"8484"
           ,x"7c04"
           ,x"0478"
           ,x"0030"
           ,x"3000"
           ,x"0030"
           ,x"3000"
           ,x"0030"
           ,x"3000"
           ,x"0030"
           ,x"1020"
           ,x"0008"
           ,x"1020"
           ,x"4020"
           ,x"1008"
           ,x"0000"
           ,x"007c"
           ,x"007c"
           ,x"0000"
           ,x"0040"
           ,x"2010"
           ,x"0810"
           ,x"2040"
           ,x"3844"
           ,x"0408"
           ,x"1010"
           ,x"0010"
           ,x"0078"
           ,x"849c"
           ,x"a498"
           ,x"807c"
           ,x"7884"
           ,x"8484"
           ,x"fc84"
           ,x"8484"
           ,x"f844"
           ,x"4478"
           ,x"4444"
           ,x"44f8"
           ,x"7884"
           ,x"8080"
           ,x"8080"
           ,x"8478"
           ,x"f844"
           ,x"4444"
           ,x"4444"
           ,x"44f8"
           ,x"fc80"
           ,x"80f0"
           ,x"8080"
           ,x"80fc"
           ,x"fc80"
           ,x"80f0"
           ,x"8080"
           ,x"8080"
           ,x"7884"
           ,x"8080"
           ,x"9c84"
           ,x"8478"
           ,x"8484"
           ,x"84fc"
           ,x"8484"
           ,x"8484"
           ,x"7c10"
           ,x"1010"
           ,x"1010"
           ,x"107c"
           ,x"0404"
           ,x"0404"
           ,x"0484"
           ,x"8478"
           ,x"8890"
           ,x"a0c0"
           ,x"a090"
           ,x"8884"
           ,x"4040"
           ,x"4040"
           ,x"4040"
           ,x"407c"
           ,x"84cc"
           ,x"b484"
           ,x"8484"
           ,x"8484"
           ,x"84c4"
           ,x"a494"
           ,x"8c84"
           ,x"8484"
           ,x"fc84"
           ,x"8484"
           ,x"8484"
           ,x"84fc"
           ,x"f884"
           ,x"8484"
           ,x"f880"
           ,x"8080"
           ,x"7884"
           ,x"8484"
           ,x"8494"
           ,x"8874"
           ,x"f884"
           ,x"8484"
           ,x"f890"
           ,x"8884"
           ,x"7884"
           ,x"8078"
           ,x"0404"
           ,x"8478"
           ,x"7c10"
           ,x"1010"
           ,x"1010"
           ,x"1010"
           ,x"8484"
           ,x"8484"
           ,x"8484"
           ,x"8478"
           ,x"4444"
           ,x"4444"
           ,x"2828"
           ,x"1010"
           ,x"8484"
           ,x"8484"
           ,x"84b4"
           ,x"cc84"
           ,x"8484"
           ,x"4830"
           ,x"3048"
           ,x"8484"
           ,x"4444"
           ,x"4428"
           ,x"1010"
           ,x"1010"
           ,x"fc04"
           ,x"0810"
           ,x"2040"
           ,x"80fc"
           ,x"3820"
           ,x"2020"
           ,x"2020"
           ,x"2038"
           ,x"0080"
           ,x"4020"
           ,x"1008"
           ,x"0400"
           ,x"7010"
           ,x"1010"
           ,x"1010"
           ,x"1070"
           ,x"1028"
           ,x"4482"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"00fc"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"544d"
           ,x"5339"
           ,x"3931"
           ,x"3035"
           ,x"2041"
           ,x"4e44"
           ,x"2046"
           ,x"5047"
           ,x"4120"
           ,x"4154"
           ,x"2057"
           ,x"4f52"
           ,x"4b21"
           ,x"2000"
           ,x"2020"
           ,x"0047"
           ,x"524f"
           ,x"4d20"
           ,x"4348"
           ,x"4543"
           ,x"4b53"
           ,x"554d"
           ,x"2054"
           ,x"4553"
           ,x"543a"
           ,x"0a0d"
           ,x"0043"
           ,x"5255"
           ,x"2046"
           ,x"524f"
           ,x"4d20"
           ,x"303a"
           ,x"2000"
           ,x"4752"
           ,x"4f4d"
           ,x"2052"
           ,x"4541"
           ,x"4420"
           ,x"5445"
           ,x"5354"
           ,x"3a31"
           ,x"3233"
           ,x"343e"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
	);
begin

	process(clk)
	variable addr_int : integer range 0 to romLast := 0;
	begin
		if rising_edge(clk) then
			addr_int := to_integer( unsigned( addr ));	-- word address
			data_out <= pgmRom( addr_int );
		end if;
	end process;

end Behavioral;
  