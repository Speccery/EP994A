----------------------------------------------------------------------------------
-- Engineer:	Erik Piehl 
-- 
-- Create Date:    07:01:30 04/15/2017 
-- Design Name: 	 testrom.vhd
-- Module Name:    testrom - Behavioral 
-- Project Name: 	 TMS9900 Test ROM code
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity testrom is
    Port ( clk : in  STD_LOGIC;
           addr : in  STD_LOGIC_VECTOR (11 downto 0);
           data_out : out  STD_LOGIC_VECTOR (15 downto 0));
end testrom;

architecture Behavioral of testrom is
	constant romLast : integer := 4095;
	type pgmRomArray is array(0 to romLast) of STD_LOGIC_VECTOR (15 downto 0);
	constant pgmRom : pgmRomArray := (  
            x"8300"
           ,x"004c"
           ,x"8380"
           ,x"0308"
           ,x"8320"
           ,x"02ca"
           ,x"beef"
           ,x"beef"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"8320"
           ,x"02f4"
           ,x"8320"
           ,x"02fe"
           ,x"0040"
           ,x"f000"
           ,x"0300"
           ,x"0002"
           ,x"020c"
           ,x"0550"
           ,x"058c"
           ,x"060c"
           ,x"0203"
           ,x"8155"
           ,x"3203"
           ,x"3603"
           ,x"0203"
           ,x"0655"
           ,x"30c3"
           ,x"04c0"
           ,x"04c1"
           ,x"0702"
           ,x"0205"
           ,x"7a9b"
           ,x"9805"
           ,x"0329"
           ,x"0204"
           ,x"000f"
           ,x"0205"
           ,x"0000"
           ,x"0206"
           ,x"f230"
           ,x"3d44"
           ,x"0204"
           ,x"000a"
           ,x"0205"
           ,x"0000"
           ,x"0206"
           ,x"0064"
           ,x"3d44"
           ,x"0206"
           ,x"0020"
           ,x"d806"
           ,x"8304"
           ,x"02ca"
           ,x"d820"
           ,x"830d"
           ,x"8305"
           ,x"02ca"
           ,x"c1e0"
           ,x"8304"
           ,x"020c"
           ,x"0400"
           ,x"04c9"
           ,x"04c2"
           ,x"d0a0"
           ,x"0324"
           ,x"0a42"
           ,x"e242"
           ,x"0b69"
           ,x"0269"
           ,x"3012"
           ,x"0202"
           ,x"0326"
           ,x"0489"
           ,x"0340"
           ,x"04c0"
           ,x"0720"
           ,x"8340"
           ,x"5820"
           ,x"031e"
           ,x"8340"
           ,x"d260"
           ,x"0320"
           ,x"1103"
           ,x"0202"
           ,x"0001"
           ,x"1001"
           ,x"0381"
           ,x"d260"
           ,x"0322"
           ,x"1101"
           ,x"10fb"
           ,x"0202"
           ,x"0011"
           ,x"0203"
           ,x"0001"
           ,x"0204"
           ,x"0002"
           ,x"3903"
           ,x"0203"
           ,x"0300"
           ,x"0204"
           ,x"5000"
           ,x"3903"
           ,x"0201"
           ,x"8000"
           ,x"0941"
           ,x"0241"
           ,x"0f00"
           ,x"0221"
           ,x"3000"
           ,x"0281"
           ,x"3a00"
           ,x"02ca"
           ,x"0201"
           ,x"b000"
           ,x"0941"
           ,x"0241"
           ,x"0f00"
           ,x"0221"
           ,x"3000"
           ,x"0281"
           ,x"3a00"
           ,x"02ca"
           ,x"0201"
           ,x"0001"
           ,x"0202"
           ,x"0002"
           ,x"8081"
           ,x"02ca"
           ,x"8042"
           ,x"02ca"
           ,x"8041"
           ,x"02ca"
           ,x"0203"
           ,x"8000"
           ,x"80c1"
           ,x"02ca"
           ,x"0704"
           ,x"80c4"
           ,x"02ca"
           ,x"c142"
           ,x"6141"
           ,x"02ca"
           ,x"c141"
           ,x"6142"
           ,x"02ca"
           ,x"c141"
           ,x"6141"
           ,x"02ca"
           ,x"0203"
           ,x"8000"
           ,x"c143"
           ,x"6141"
           ,x"02ca"
           ,x"0704"
           ,x"c143"
           ,x"6144"
           ,x"02ca"
           ,x"0420"
           ,x"0008"
           ,x"020c"
           ,x"0240"
           ,x"1d00"
           ,x"0202"
           ,x"0001"
           ,x"288c"
           ,x"20a0"
           ,x"0048"
           ,x"1301"
           ,x"0381"
           ,x"24a0"
           ,x"004a"
           ,x"1301"
           ,x"0381"
           ,x"1d00"
           ,x"1e01"
           ,x"1d02"
           ,x"1eff"
           ,x"1f00"
           ,x"1301"
           ,x"0381"
           ,x"1f01"
           ,x"1601"
           ,x"0381"
           ,x"0200"
           ,x"3333"
           ,x"2c20"
           ,x"beef"
           ,x"0200"
           ,x"5555"
           ,x"2c60"
           ,x"0011"
           ,x"020c"
           ,x"0550"
           ,x"0203"
           ,x"0055"
           ,x"3003"
           ,x"3243"
           ,x"0203"
           ,x"0006"
           ,x"0a83"
           ,x"30c3"
           ,x"04cc"
           ,x"0208"
           ,x"0012"
           ,x"3608"
           ,x"3409"
           ,x"0288"
           ,x"7912"
           ,x"1301"
           ,x"0381"
           ,x"0289"
           ,x"a079"
           ,x"1301"
           ,x"0381"
           ,x"0203"
           ,x"8340"
           ,x"0207"
           ,x"8350"
           ,x"0201"
           ,x"0123"
           ,x"0202"
           ,x"4567"
           ,x"0204"
           ,x"89ab"
           ,x"c4c1"
           ,x"c8c2"
           ,x"0002"
           ,x"c8c4"
           ,x"0004"
           ,x"04e3"
           ,x"0006"
           ,x"ddf3"
           ,x"ddf3"
           ,x"ddf3"
           ,x"ddf3"
           ,x"cdf3"
           ,x"d820"
           ,x"8303"
           ,x"8350"
           ,x"0203"
           ,x"8340"
           ,x"d804"
           ,x"8340"
           ,x"d802"
           ,x"8341"
           ,x"c4c1"
           ,x"d4c4"
           ,x"bcc1"
           ,x"b4c1"
           ,x"0223"
           ,x"ffff"
           ,x"d073"
           ,x"d053"
           ,x"0603"
           ,x"04d3"
           ,x"0204"
           ,x"8350"
           ,x"0202"
           ,x"0002"
           ,x"cd33"
           ,x"0644"
           ,x"ad02"
           ,x"6802"
           ,x"8350"
           ,x"0283"
           ,x"8342"
           ,x"1301"
           ,x"0381"
           ,x"0201"
           ,x"4444"
           ,x"c801"
           ,x"8360"
           ,x"c820"
           ,x"8360"
           ,x"8350"
           ,x"8060"
           ,x"8350"
           ,x"1301"
           ,x"0381"
           ,x"0200"
           ,x"1234"
           ,x"0381"
           ,x"06a0"
           ,x"02c4"
           ,x"04c1"
           ,x"04e3"
           ,x"0004"
           ,x"0723"
           ,x"0006"
           ,x"04e0"
           ,x"8348"
           ,x"0713"
           ,x"04f3"
           ,x"04f3"
           ,x"04f3"
           ,x"0502"
           ,x"ccc2"
           ,x"10f0"
           ,x"0502"
           ,x"0202"
           ,x"8002"
           ,x"0502"
           ,x"0502"
           ,x"05c3"
           ,x"c143"
           ,x"0585"
           ,x"0605"
           ,x"06c5"
           ,x"0545"
           ,x"0713"
           ,x"0745"
           ,x"0505"
           ,x"0200"
           ,x"1234"
           ,x"0201"
           ,x"0001"
           ,x"c4c0"
           ,x"c0b3"
           ,x"a081"
           ,x"c202"
           ,x"c4c1"
           ,x"a4c1"
           ,x"c820"
           ,x"0004"
           ,x"8344"
           ,x"06a0"
           ,x"02c4"
           ,x"0460"
           ,x"004c"
           ,x"0204"
           ,x"007b"
           ,x"045b"
           ,x"03a0"
           ,x"02a0"
           ,x"0202"
           ,x"0004"
           ,x"c0c2"
           ,x"0583"
           ,x"6083"
           ,x"02c1"
           ,x"0200"
           ,x"0004"
           ,x"c040"
           ,x"0202"
           ,x"fffc"
           ,x"c0c0"
           ,x"0204"
           ,x"fffc"
           ,x"0a81"
           ,x"0812"
           ,x"0b43"
           ,x"0914"
           ,x"0380"
           ,x"020c"
           ,x"0100"
           ,x"02c1"
           ,x"1d00"
           ,x"0380"
           ,x"020c"
           ,x"0100"
           ,x"02c1"
           ,x"1d01"
           ,x"0380"
           ,x"0200"
           ,x"4455"
           ,x"0201"
           ,x"6677"
           ,x"02ca"
           ,x"0380"
           ,x"d040"
           ,x"02ca"
           ,x"d080"
           ,x"02ca"
           ,x"045b"
           ,x"2080"
           ,x"4000"
           ,x"a000"
           ,x"0800"
           ,x"0c00"
           ,x"8090"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
           ,x"0000"
	);
begin

	process(clk)
	variable addr_int : integer range 0 to romLast := 0;
	begin
		if rising_edge(clk) then
			addr_int := to_integer( unsigned( addr ));	-- word address
			data_out <= pgmRom( addr_int );
		end if;
	end process;

end Behavioral;
  